module translator_update (
        input  logic        i_clk, i_reset,
        input  logic [15:0] i_toDisplay_bin,
        output logic        o_update
    );

    logic [15:0] pr_input, nx_input;

    

endmodule;