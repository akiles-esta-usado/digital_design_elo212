`timescale 1ns / 1ps

module tb_top_2 ();

endmodule