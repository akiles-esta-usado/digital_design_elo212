`timescale 1ns / 1ps

module S4_Actividad3 (

);
    
endmodule