`timescale 1ns / 1ps

module semaforoTimer #(parameter DELAY = 5) (
	input  logic       clock,
	input  logic       reset, TA, TB,
	output logic [1:0] LA, LB);

    localparam DELAY_WIDTH = $clog2(DELAY);
	logic [DELAY_WIDTH-1:0]  delay_timer;
	
    enum logic[3:0] {
        STATE_0 = 4'b0001,
        STATE_1 = 4'b0010,
        STATE_2 = 4'b0100,
        STATE_3 = 4'b1000
        } state, next_state;
    
    //output encoding
    localparam GREEN    = 2'b00;
    localparam YELLOW   = 2'b01;
    localparam RED      = 2'b10;
    
    always_ff @(posedge clock) begin
        if (reset) delay_timer <= 0;
        else if (state != next_state) delay_timer <= 0; // reset the timer when state changes
        else delay_timer <= delay_timer + 1;
    end
    
    // one combinational block computes the next_state and outputs for the
    // current state
    always_comb begin
        //using default assignments here allows us to save space, helps on readability,
        //and reduces the chance of unintentional errors
        next_state = state;
    	LA = RED;
    	LB = RED;
    	
    	case (state)
    		STATE_0: begin
    			     LA = GREEN;
    			     if(TA == 1'b0 && (delay_timer >= DELAY-1)) begin
    			 	   next_state = STATE_1;
    		         end
    		    end

            STATE_1: begin
                    LA = YELLOW;
                    if(delay_timer >= DELAY-1) begin
    			 	   next_state = STATE_2;
    		        end

                end
            
            STATE_2: begin
                    LB = GREEN;
                    if(TB == 1'b0 && (delay_timer >= DELAY-1)) begin
                        next_state = STATE_3;
                    end
                end

            STATE_3: begin
                    LB = YELLOW;
                    if(delay_timer >= DELAY-1) begin
    			 	   next_state = STATE_0;
    		        end
                end                
    	endcase
    end	

    // when clock ticks, update the state
    always_ff @(posedge clock) begin
    	if(reset) state <= STATE_0;
    	else state <= next_state;
    end
endmodule