`timescale 1ns / 1ps

module tb_mux_4(

    );
endmodule
