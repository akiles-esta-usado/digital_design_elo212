`timescale 1ns / 1ps

module tb_top_3 ();

endmodule