`timescale 1ns / 1ps

module tb_top_1 ();

endmodule