`timescale 1ns / 1ps



module tb_new_testbench();

    logic clk, reset;

    // 
    logic in, out;

endmodule


module reader(
        input  logic i_clk, i_reset;
        input  logic i_in;
        output logic o_out;
        );


endmodule


module signal_generator(
        input  logic i_clk, i_reset;
        );


endmodule


module verifier(
        input  logic i_clk, i_reset;
        input  logic   in;
        );

endmodule
